module Lab2_4_bit_BLS_dataflow(input [3:0] A,B, input bin, output [3:0] D, output bout);
    assign D[0] = (A[0])^(B[0])^(bin),
           D[1] = (A[1])^(B[1])^((~(A[0]^B[0])&bin)|((~A[0])&B[0])),
           D[2] = (A[2])^(B[2])^(((~(A[1]^B[1])&((~(A[0]^B[0])&bin)|((~A[0])&B[0])))|((~A[1])&B[1]))),
           D[3] = (A[3])^(B[3])^(((~(A[2]^B[2])&(((~(A[1]^B[1])&((~(A[0]^B[0])&bin)|((~A[0])&B[0])))|((~A[1])&B[1]))))|((~A[2])&B[2]))),

           bout = ((~(A[3]^B[3])&(((~(A[2]^B[2])&(((~(A[1]^B[1])&((~(A[0]^B[0])&bin)|((~A[0])&B[0])))|((~A[1])&B[1]))))|((~A[2])&B[2]))))|((~A[3])&B[3]));

endmodule

        //    b0 = bin
        //    b1 = ((~(A[0]^B[0])&bin)|((~A[0])&B[0]))
        //    b2 = (((~(A[1]^B[1])&((~(A[0]^B[0])&bin)|((~A[0])&B[0])))|((~A[1])&B[1])))
        //    b3 = (((~(A[2]^B[2])&(((~(A[1]^B[1])&((~(A[0]^B[0])&bin)|((~A[0])&B[0])))|((~A[1])&B[1]))))|((~A[2])&B[2])))

module Lab1_gatelevel_UDP(F,A,B,C,D);
    output  F;
    input   A,B,C,D;

    Lab1_UDP M0(F,A,B,C,D);


endmodule